// to use insAI extension
`define ENABLE_insAI_EXTENSION 
